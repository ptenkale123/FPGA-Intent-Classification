module testbench();

timeunit 10ns;	

timeprecision 1ns;

logic in;
logic out;
nn_wrapper dut (.*);

endmodule
