nn_partition p_1 (.*,
.W_1(32'hbe0b7026), .W_2(32'hbdf58e22), .W_3(32'hbd857215), .W_4(32'hbdd2ec6c), 
.W_5(32'h3c223183), .W_6(32'h3d98d930), .W_7(32'hbb098f60), .W_8(32'h3cf9ce8e), 
.W_9(32'hbd967fd4), .W_10(32'h3d848494), .W_11(32'h3c06ab80), .W_12(32'h3ce9984a), 
.W_13(32'h3c52b2c0), .W_14(32'h3ccc5543), .W_15(32'h3c03b4c0), .W_16(32'h3e0a6a01), 
.W_17(32'hbd2bde40), .W_18(32'h3d23c85c), .W_19(32'h3da24fec), .W_20(32'hbd8d7492), 
.W_21(32'hbcad8c2a), .W_22(32'h3bc58256), .W_23(32'h3c0c8abd), .W_24(32'h3d37c569), 
.W_25(32'h3c0bc7b4), .W_26(32'hbd856cd7), .W_27(32'h3cd245b3), .W_28(32'hbddefc7a), 
.W_29(32'h3bf3ee7a), .W_30(32'hbd84aa54), .W_31(32'h3d284381), .W_32(32'h3d5947d0), 
.W_33(32'h3d76848c), .W_34(32'hbd8ffb8b), .W_35(32'hbcb01c93), .W_36(32'hbc0ba4e4), 
.W_37(32'hbc733440), .W_38(32'h3cbeec39), .W_39(32'hbd15feda), .W_40(32'h3c670c13), 
.W_41(32'hbcdeedcc), .W_42(32'hbd8e4b02), .W_43(32'hbcb1012a), .W_44(32'hbe06f156), 
.W_45(32'h3da3aeab), .W_46(32'h3d80a5ad), .W_47(32'h3d81986c), .W_48(32'hbdae4218), 
.W_49(32'hbc1c220a), .W_50(32'hbc8be511), .W_51(32'hbd9d04a3), .W_52(32'hbd874ea9), 
.W_53(32'h3d65adda), .W_54(32'hbdbd6b66), .W_55(32'h3d3892ef), .W_56(32'hbd2b4c7f), 
.W_57(32'hbd39da16), .W_58(32'hbde9003f), .W_59(32'h3d0e3bcd), .W_60(32'hbd8846a6), 
.W_61(32'h3d7d5886), .W_62(32'hbdd2f6e8), .W_63(32'hbddddc1e), .W_64(32'hbd1aee63), 
.bias(32'hbe4cb296), .out(O_1));

nn_partition p_2 (.*,
.W_1(32'hbe4cba73), .W_2(32'hbc6f5233), .W_3(32'h3c113cd4), .W_4(32'h3ca8ae75), 
.W_5(32'hbeaf583a), .W_6(32'hbdcd844d), .W_7(32'h3e06833c), .W_8(32'hbdf1bef5), 
.W_9(32'hbdfdb4cc), .W_10(32'hbbe14021), .W_11(32'h3c1e0462), .W_12(32'h3d4621b8), 
.W_13(32'h3d2310dc), .W_14(32'h3cc3f5f9), .W_15(32'h3b6cad3d), .W_16(32'h3cae48e9), 
.W_17(32'h3c56cb53), .W_18(32'hbd94256c), .W_19(32'hbd013fd1), .W_20(32'hbccb599b), 
.W_21(32'hbda6aa8f), .W_22(32'h3d02cd3a), .W_23(32'hbc5527e5), .W_24(32'h3ce4bec6), 
.W_25(32'hbd03b2dd), .W_26(32'hbd68ef78), .W_27(32'h3d8408d9), .W_28(32'h3c1e4b45), 
.W_29(32'hbd33b646), .W_30(32'hbdc90710), .W_31(32'hbc979182), .W_32(32'h3cdbab22), 
.W_33(32'hbc57f51f), .W_34(32'h3d0d0cc3), .W_35(32'hbb997ec2), .W_36(32'hbd020e63), 
.W_37(32'hbdcab713), .W_38(32'h3d28c693), .W_39(32'h3d3152f4), .W_40(32'hbd88c500), 
.W_41(32'h3d3f3e03), .W_42(32'hbd91e8e6), .W_43(32'hbd135547), .W_44(32'hbd9bccaf), 
.W_45(32'hbc52d44e), .W_46(32'hbc920e1f), .W_47(32'h3c4bd556), .W_48(32'hbd2c28b3), 
.W_49(32'hbdaf5d35), .W_50(32'hbbf32f37), .W_51(32'h3c988b11), .W_52(32'h3db7c569), 
.W_53(32'h3d5691a7), .W_54(32'hbdbb00bd), .W_55(32'hbc91fb40), .W_56(32'h3c39f55a), 
.W_57(32'hbd77a3db), .W_58(32'hbe18ab0d), .W_59(32'hbd16cb53), .W_60(32'h3ce9d94d), 
.W_61(32'hbd993ee6), .W_62(32'hbd64b33e), .W_63(32'hbda29739), .W_64(32'hbd42e01a), 
.bias(32'hbf1b22d1), .out(O_2));

nn_partition p_3 (.*,
.W_1(32'h3d944f5d), .W_2(32'hbdbfb2ee), .W_3(32'hbd540358), .W_4(32'hbe1923a3), 
.W_5(32'h3d4d0edc), .W_6(32'h3c3acb43), .W_7(32'hbbbc6145), .W_8(32'h3c6425af), 
.W_9(32'h3ceeb0b8), .W_10(32'h3d112dba), .W_11(32'h3cc92360), .W_12(32'h3d8343b7), 
.W_13(32'h3c9d4952), .W_14(32'h3dcece9a), .W_15(32'h3d6b6ae8), .W_16(32'h3ca0e842), 
.W_17(32'h3bbc2911), .W_18(32'hbb1e5413), .W_19(32'h3daea20a), .W_20(32'h3ce9b38d), 
.W_21(32'hbc39d3cc), .W_22(32'hbc70f16f), .W_23(32'h3d43ad9f), .W_24(32'h3d415a08), 
.W_25(32'h3c82517e), .W_26(32'hbb976435), .W_27(32'h3dc4e1e7), .W_28(32'hbd317375), 
.W_29(32'h3dedea89), .W_30(32'hbac3b0c4), .W_31(32'h3ce11340), .W_32(32'h3db7f280), 
.W_33(32'h3d458dde), .W_34(32'hbd3c2fc7), .W_35(32'hbd7d4e09), .W_36(32'h3cbd640f), 
.W_37(32'hb7a9f850), .W_38(32'h3d72cd7d), .W_39(32'h3cd4690e), .W_40(32'h3af1a198), 
.W_41(32'h3d36c69b), .W_42(32'hbd4e4a7b), .W_43(32'hbd6a64c3), .W_44(32'hbd79f87f), 
.W_45(32'h3d357a35), .W_46(32'hbb3266f0), .W_47(32'h3dccb641), .W_48(32'h3c4d6c2f), 
.W_49(32'hbc2a1512), .W_50(32'h3c72d3c8), .W_51(32'h3d2cd5b7), .W_52(32'h3d7264a1), 
.W_53(32'h3cedf1e1), .W_54(32'hbdc1b64e), .W_55(32'h3df89614), .W_56(32'hbcb2f230), 
.W_57(32'h3d0f41f2), .W_58(32'hbd606a6e), .W_59(32'h3e16555c), .W_60(32'h3d90afe6), 
.W_61(32'h3dade764), .W_62(32'h398f59d0), .W_63(32'h3d417b96), .W_64(32'h4012b1c4), 
.bias(32'h3ef60419), .out(O_3));

