nn_partition p_1 (.*,
.W_1(32'h3f588e37), .W_2(32'hbd106141), .W_3(32'hbd1a0275), .W_4(32'hbd3a0a52), 
.W_5(32'h3e17bf1f), .W_6(32'h3c82b40f), .W_7(32'h3e06defc), .W_8(32'h3dfc4b0a), 
.W_9(32'hbe37342f), .W_10(32'hbdb2b021), .W_11(32'hbdbe5754), .W_12(32'hbcebf013), 
.W_13(32'hbdb1c53f), .W_14(32'h3d965a9b), .W_15(32'hbe375643), .W_16(32'hbe41450f), 
.W_17(32'h3bc9978e), .W_18(32'hbdb91a33), .W_19(32'hbe094706), .W_20(32'hbd9f394b), 
.W_21(32'hbe089ca2), .W_22(32'hbc643244), .W_23(32'hbdf404ea), .W_24(32'hbda59ea5), 
.W_25(32'hbda9a4df), .W_26(32'hbdbcd0bb), .W_27(32'hbe02db62), .W_28(32'hbd2ab25b), 
.W_29(32'hbd3a82e8), .W_30(32'hbd10ecb7), .W_31(32'hbdb4213a), .W_32(32'hbdac35ce), 
.W_33(32'hbd6733ec), .W_34(32'hbd9a4053), .W_35(32'hbe0c2507), .W_36(32'hbd7be985), 
.W_37(32'hbdb821af), .W_38(32'hbd7fc548), .W_39(32'hbcfe1544), .W_40(32'hbd203d57), 
.W_41(32'hbd21e929), .W_42(32'hbd8c2374), .W_43(32'hbd064ba9), .W_44(32'hbd00c73b), 
.W_45(32'hbd0d79d1), .W_46(32'h3c0701e7), .W_47(32'hbd9a4378), .W_48(32'hbd71d92b), 
.W_49(32'hbd95e072), .W_50(32'hbdb2684d), .W_51(32'hbdc99ae9), .W_52(32'h3bedc139), 
.W_53(32'hbd812d77), .W_54(32'h3a7ef6c1), .W_55(32'hbd289225), .W_56(32'h3c6cd4aa), 
.W_57(32'h3d8bf4cb), .W_58(32'h3c923e5c), .W_59(32'h3ce2f9ca), .W_60(32'hbd09ce4a), 
.W_61(32'h3d3fdb4d), .W_62(32'h3dba786c), .W_63(32'hbb9b0ee5), .W_64(32'h3d0ee8d1), 
.bias(32'h3f55f6fd), .out(O_1));

nn_partition p_2 (.*,
.W_1(32'hbf26ee0f), .W_2(32'h3db5dcc6), .W_3(32'h3ef4816f), .W_4(32'h3ed0f51b), 
.W_5(32'h3a1b9e82), .W_6(32'h3e679bbb), .W_7(32'hbe505293), .W_8(32'hbe88d3ae), 
.W_9(32'h3c203a32), .W_10(32'hbea6f156), .W_11(32'h3ea8754f), .W_12(32'hbcfca85d), 
.W_13(32'hbd170d63), .W_14(32'hbdb1b2e6), .W_15(32'h3e45ac47), .W_16(32'h3e8b2570), 
.W_17(32'h3d708787), .W_18(32'h3df8ca82), .W_19(32'h3d45e6ff), .W_20(32'h3d337111), 
.W_21(32'h3e44e50c), .W_22(32'h3d80181e), .W_23(32'hbe0f27bb), .W_24(32'h3e875a32), 
.W_25(32'h3da33a47), .W_26(32'h3e0877ee), .W_27(32'h3d90aaa8), .W_28(32'h3e5458cd), 
.W_29(32'h3e2bde40), .W_30(32'h3df75105), .W_31(32'h3dbd6a59), .W_32(32'h3e80e022), 
.W_33(32'h3d1f3e8a), .W_34(32'hbd691ea8), .W_35(32'h3e287fcc), .W_36(32'hbe4548aa), 
.W_37(32'h3ddba0a5), .W_38(32'hbdb0d38d), .W_39(32'hbdce703b), .W_40(32'hbd333b97), 
.W_41(32'h3d8ea077), .W_42(32'hbd85870e), .W_43(32'hbe79652c), .W_44(32'hbdcb3dd1), 
.W_45(32'h3dd3cddd), .W_46(32'hbd09c2c2), .W_47(32'hbe11af3a), .W_48(32'hbcd000c9), 
.W_49(32'h3d82e01a), .W_50(32'hbc74adbc), .W_51(32'hbd58d8a9), .W_52(32'h3da5c897), 
.W_53(32'hbe027d03), .W_54(32'hbdd7396d), .W_55(32'h3dab4e12), .W_56(32'hbd3865d8), 
.W_57(32'hbe40c49c), .W_58(32'hbdf8476f), .W_59(32'hbe7ce853), .W_60(32'h3d704791), 
.W_61(32'hbe6e410b), .W_62(32'hbd3c45cc), .W_63(32'hbe1b90eb), .W_64(32'hbe8415f4), 
.bias(32'hbf085879), .out(O_2));

nn_partition p_3 (.*,
.W_1(32'h3e77e3d2), .W_2(32'h3d3aa79c), .W_3(32'hbe35da27), .W_4(32'hbe3559b4), 
.W_5(32'h3d81fc8f), .W_6(32'hbdc1b973), .W_7(32'h3e8342ee), .W_8(32'h3eacbe62), 
.W_9(32'h3e55feda), .W_10(32'h3dac4bd3), .W_11(32'hbe31f362), .W_12(32'h3f1b7d41), 
.W_13(32'h3eaa2f06), .W_14(32'h3e3a1230), .W_15(32'h3e0eac86), .W_16(32'h3e4a4a8c), 
.W_17(32'h3e530404), .W_18(32'h3ecb9b67), .W_19(32'h3ec44d01), .W_20(32'h3e43a53c), 
.W_21(32'h3e06fe72), .W_22(32'h3e3fb15b), .W_23(32'h3ea83904), .W_24(32'h3e6f227d), 
.W_25(32'h3ea80dc3), .W_26(32'h3e1ebaf1), .W_27(32'h3e0dc875), .W_28(32'h3dc86727), 
.W_29(32'h3e19abf3), .W_30(32'h3e1e132b), .W_31(32'h3e489763), .W_32(32'h3e234eba), 
.W_33(32'h3e3ab9f5), .W_34(32'h3d05b39e), .W_35(32'h3e1cb3e5), .W_36(32'h3ce47bab), 
.W_37(32'h3cd95bbc), .W_38(32'hbc2d6883), .W_39(32'hbd456606), .W_40(32'hbd68b5cc), 
.W_41(32'hbde339c1), .W_42(32'hbce2e903), .W_43(32'hbcdf82b2), .W_44(32'hbd8abf77), 
.W_45(32'hbdc3d4f1), .W_46(32'hbdb39757), .W_47(32'h3b6ebdb8), .W_48(32'hbe01d53d), 
.W_49(32'h39893777), .W_50(32'hbdf15619), .W_51(32'hbd87b4e5), .W_52(32'hbd8d1b71), 
.W_53(32'hbcbcf701), .W_54(32'hbdf266ba), .W_55(32'hbe1bdcf0), .W_56(32'hbdaa4b99), 
.W_57(32'h3d9f79c8), .W_58(32'h3d18d691), .W_59(32'h3ca8e2e3), .W_60(32'hbe0bce85), 
.W_61(32'h3bbd8531), .W_62(32'hbd8daa0d), .W_63(32'h3d92a066), .W_64(32'h3de7b0b4), 
.bias(32'h3d99ce07), .out(O_3));

nn_partition p_4 (.*,
.W_1(32'hbf0b0be1), .W_2(32'hbdcb0c89), .W_3(32'h3e372c52), .W_4(32'h3de6d9be), 
.W_5(32'hbdedefc8), .W_6(32'h3de415f4), .W_7(32'hbe866517), .W_8(32'hbe9ca81a), 
.W_9(32'hbe56bb99), .W_10(32'hbe36fd22), .W_11(32'h3f2f1d3f), .W_12(32'h3e8d844d), 
.W_13(32'h3e8ac322), .W_14(32'h3d857753), .W_15(32'h3e86b26c), .W_16(32'hbea3a7db), 
.W_17(32'h3b0ae8fd), .W_18(32'h3e7f9f02), .W_19(32'h3d52274a), .W_20(32'hbda54ac3), 
.W_21(32'h3d4d2d45), .W_22(32'h3d68fe26), .W_23(32'h3dc5e3da), .W_24(32'hbcfb9e06), 
.W_25(32'h3e52a844), .W_26(32'h3e13a14d), .W_27(32'h3ece108c), .W_28(32'h3e5bbadc), 
.W_29(32'h3e1ce315), .W_30(32'h3da9a134), .W_31(32'h3e929b28), .W_32(32'hbd8594af), 
.W_33(32'h3e15e204), .W_34(32'h3d631833), .W_35(32'hbb869d3e), .W_36(32'h3e28a71e), 
.W_37(32'h3e09613d), .W_38(32'h3d054ef4), .W_39(32'h3de45f5b), .W_40(32'h3d2aa194), 
.W_41(32'hbdf68f08), .W_42(32'h3e2995ab), .W_43(32'hbd6379b7), .W_44(32'h3da699c8), 
.W_45(32'h3d966cf4), .W_46(32'h3da345d0), .W_47(32'hbd868a93), .W_48(32'h3e427fa2), 
.W_49(32'hbba5947a), .W_50(32'h3d7abda1), .W_51(32'hbe1bf488), .W_52(32'hbdb3061c), 
.W_53(32'h3df47d80), .W_54(32'h3dd2934b), .W_55(32'hbd0e8b7e), .W_56(32'h3cc93a71), 
.W_57(32'h3c021ebe), .W_58(32'h3dc82f94), .W_59(32'hbe21cac1), .W_60(32'hbe75c7ce), 
.W_61(32'hbc62c55d), .W_62(32'h3e107f24), .W_63(32'hbd6188b1), .W_64(32'hbd0a01ac), 
.bias(32'hbf24c986), .out(O_4));

nn_partition p_5 (.*,
.W_1(32'hbf32dcb1), .W_2(32'h3d3e4ef0), .W_3(32'h3eae410b), .W_4(32'h3e8f1bef), 
.W_5(32'h3cac710d), .W_6(32'hbe0b4396), .W_7(32'hbd1ba5e3), .W_8(32'hbcfea3df), 
.W_9(32'hbe4afa2f), .W_10(32'hbd7074a7), .W_11(32'h3d87b4e5), .W_12(32'hbddeb852), 
.W_13(32'h3d3b7e91), .W_14(32'hbeafe9b8), .W_15(32'hbeae8d11), .W_16(32'hbe5d1245), 
.W_17(32'hbec400fc), .W_18(32'hbe85c52e), .W_19(32'hbefa3593), .W_20(32'hbee7136a), 
.W_21(32'hbeba0126), .W_22(32'hbed0e172), .W_23(32'hbe64c597), .W_24(32'hbed58256), 
.W_25(32'hbeb5158c), .W_26(32'hbe9cd9e8), .W_27(32'hbef04ab6), .W_28(32'hbe702de0), 
.W_29(32'hbf11aaa4), .W_30(32'hbe9e69ad), .W_31(32'hbeb17ebb), .W_32(32'hbe91d53d), 
.W_33(32'hbec22920), .W_34(32'hbe57e133), .W_35(32'hbe29fbe7), .W_36(32'hbdd374bc), 
.W_37(32'hbc8ed1bf), .W_38(32'h3cc9949f), .W_39(32'h3ca0663c), .W_40(32'h3d450df1), 
.W_41(32'h3e1fa440), .W_42(32'h3a7a8699), .W_43(32'hbd8bb342), .W_44(32'h3d32ebe6), 
.W_45(32'h3d509e13), .W_46(32'h3be7eb36), .W_47(32'h3b26f09a), .W_48(32'hbd4bcf0b), 
.W_49(32'hbc01b7fc), .W_50(32'hbbfb3df9), .W_51(32'h3cae2fbe), .W_52(32'h3d3394b8), 
.W_53(32'hbdd58b82), .W_54(32'h3c62046c), .W_55(32'h3cb73d19), .W_56(32'h3d786a0a), 
.W_57(32'h3d0fcb4f), .W_58(32'hbcf7dfa0), .W_59(32'h3cef501a), .W_60(32'hbcd71d1d), 
.W_61(32'h3dc0a5ad), .W_62(32'h3dbb267c), .W_63(32'hbd904e62), .W_64(32'hbc0544e3), 
.bias(32'hbf3ccccd), .out(O_5));

nn_partition p_6 (.*,
.W_1(32'hbece2047), .W_2(32'h3deeb702), .W_3(32'hbe383516), .W_4(32'hbdea5508), 
.W_5(32'h3d61198b), .W_6(32'h3db15f89), .W_7(32'h3f2c6888), .W_8(32'hbe991fb4), 
.W_9(32'h3d676b7f), .W_10(32'hbe941355), .W_11(32'hbf03b44e), .W_12(32'hbed0370d), 
.W_13(32'hbe98d10f), .W_14(32'hbd40431c), .W_15(32'h3e99a954), .W_16(32'h3eba2c67), 
.W_17(32'h3e923e18), .W_18(32'hbe22aed1), .W_19(32'h3d82cc2d), .W_20(32'h3e7436b9), 
.W_21(32'h3e7cbe62), .W_22(32'h3ea9e98e), .W_23(32'hbda3b57c), .W_24(32'h3e13bb84), 
.W_25(32'h3d0da3c2), .W_26(32'hbdc1c609), .W_27(32'hbe06277c), .W_28(32'h3d87032a), 
.W_29(32'h3d6b4fa5), .W_30(32'h3e7fa97e), .W_31(32'h3e6ba1f5), .W_32(32'hbcd0c804), 
.W_33(32'hbd8240b8), .W_34(32'hbc35cbff), .W_35(32'hbcc97b74), .W_36(32'h3e23b795), 
.W_37(32'h3e208d8f), .W_38(32'h3e3f4342), .W_39(32'h3e18ab0d), .W_40(32'hbd31b047), 
.W_41(32'h3d872431), .W_42(32'hbcd8adac), .W_43(32'hbd262cba), .W_44(32'hbc22edd6), 
.W_45(32'h3d209dd0), .W_46(32'h3c0cd856), .W_47(32'h3cddd2af), .W_48(32'hbdef1aa0), 
.W_49(32'h3e705293), .W_50(32'h3e4493c9), .W_51(32'h3d94a904), .W_52(32'hbd5e3865), 
.W_53(32'h3e355c53), .W_54(32'h3cd985ad), .W_55(32'h3ae8ed95), .W_56(32'h3e3f62b7), 
.W_57(32'h3da941c8), .W_58(32'hbdf5d24a), .W_59(32'h3e22602d), .W_60(32'hbd3d9a95), 
.W_61(32'h3e84894c), .W_62(32'h3dcc94b4), .W_63(32'hbd762952), .W_64(32'h3e045cbc), 
.bias(32'hbe31de6a), .out(O_6));

nn_partition p_7 (.*,
.W_1(32'hbf680735), .W_2(32'hbe2b09ea), .W_3(32'h3e83d5bb), .W_4(32'h3f2e108c), 
.W_5(32'hbe33ae68), .W_6(32'h3da5da6a), .W_7(32'hbe0b5b2d), .W_8(32'hbd167664), 
.W_9(32'h3f47c06e), .W_10(32'h3e2beb5b), .W_11(32'h3f54da90), .W_12(32'h3e804ff4), 
.W_13(32'h3e2255b0), .W_14(32'h3ddd0a67), .W_15(32'h3ecf598a), .W_16(32'h3ea82a99), 
.W_17(32'hbcdc7043), .W_18(32'h3e4b9cb7), .W_19(32'h3e073ffb), .W_20(32'h3be708b8), 
.W_21(32'h3ef599ed), .W_22(32'hb9414606), .W_23(32'h3e113be2), .W_24(32'h3e8f9485), 
.W_25(32'h3edfa58f), .W_26(32'h3e9039ac), .W_27(32'h3d1c054f), .W_28(32'h3e98ac5c), 
.W_29(32'h3e4400fc), .W_30(32'h3e931ceb), .W_31(32'h3f21de6a), .W_32(32'h3e492253), 
.W_33(32'h3e9cf41f), .W_34(32'h3ea5d639), .W_35(32'h3d085d31), .W_36(32'h3f00793e), 
.W_37(32'h3eb30942), .W_38(32'h3c9374bc), .W_39(32'h3e783cf3), .W_40(32'h3e9b83cf), 
.W_41(32'h3edede55), .W_42(32'h3ea47065), .W_43(32'h3ed1719f), .W_44(32'h3e939970), 
.W_45(32'h3e41e4f7), .W_46(32'h3e39c38b), .W_47(32'h3ebcd4aa), .W_48(32'h3e85fd8b), 
.W_49(32'h3e71fddf), .W_50(32'h3e213554), .W_51(32'h3e64ab60), .W_52(32'h3ed1758e), 
.W_53(32'h3e0aa8eb), .W_54(32'h3db3ade2), .W_55(32'h3d033e79), .W_56(32'h3e8d7c70), 
.W_57(32'h3e4c5eb3), .W_58(32'h3de6eeb7), .W_59(32'h3e3d5bab), .W_60(32'h3d862802), 
.W_61(32'h3e97e282), .W_62(32'h3e37d6b6), .W_63(32'h3e3e83e4), .W_64(32'h3e605921), 
.bias(32'hbf3b4396), .out(O_7));

nn_partition p_8 (.*,
.W_1(32'hbf72599f), .W_2(32'h3f4fe719), .W_3(32'hbe1f40a3), .W_4(32'hbe052e73), 
.W_5(32'h3f5d551d), .W_6(32'hbe9f05a7), .W_7(32'h3ec8d64d), .W_8(32'hbf691d15), 
.W_9(32'h3cac2bd8), .W_10(32'h3f5760bf), .W_11(32'h3da9c348), .W_12(32'hbe4dbb5a), 
.W_13(32'hbf0db61c), .W_14(32'hbe861523), .W_15(32'hbdcbf3bf), .W_16(32'h3e5251c2), 
.W_17(32'h3e4caff7), .W_18(32'h3e39a416), .W_19(32'hbd1287c2), .W_20(32'h3ec0a527), 
.W_21(32'h3eed7881), .W_22(32'h3e50ff97), .W_23(32'h3e07381d), .W_24(32'h3df73190), 
.W_25(32'h3e195033), .W_26(32'h3df7fe09), .W_27(32'hbd29ec2d), .W_28(32'hbcdd4e90), 
.W_29(32'hbdfc6a7f), .W_30(32'h3d2fcdee), .W_31(32'h3d902603), .W_32(32'h3e0e7818), 
.W_33(32'h3df290ac), .W_34(32'h3e89081c), .W_35(32'h3e23a53c), .W_36(32'h3db02e66), 
.W_37(32'h3b022e43), .W_38(32'hbd5ca6ca), .W_39(32'h3e21205c), .W_40(32'h3d48c826), 
.W_41(32'h3e086595), .W_42(32'hbdb6cc60), .W_43(32'h3dcc6de7), .W_44(32'hbd8b4528), 
.W_45(32'h3d50b73d), .W_46(32'h3dcea9e7), .W_47(32'h3e299d88), .W_48(32'hbe3d70a4), 
.W_49(32'h3e225aee), .W_50(32'h3dbb9f99), .W_51(32'h3da91fb4), .W_52(32'h3dff62b7), 
.W_53(32'hbd5f6662), .W_54(32'h3d44816f), .W_55(32'h3e9754f3), .W_56(32'h3d279fed), 
.W_57(32'hbe08f323), .W_58(32'hbdade43f), .W_59(32'h3e5b6c37), .W_60(32'h3dba005c), 
.W_61(32'h3cca6ca0), .W_62(32'h3dc4a9ce), .W_63(32'hbd05cee1), .W_64(32'hbd5c7ef1), 
.bias(32'hbf48240b), .out(O_8));

